`timescale 1ns/100ps

module Array_44 #(
	parameter DATA_WIDTH = 8,
	parameter BLOCK_SIZE = 4,
	parameter SELECT_WIDTH = 2,
	parameter ARRAY_SIZE = 4
	)(
	input [BLOCK_SIZE*BLOCK_SIZE*DATA_WIDTH-1:0]Input_act[ARRAY_SIZE-1:0],
	input [DATA_WIDTH-1:0]Input_weight[ARRAY_SIZE-1:0],
	input [DATA_WIDTH-1:0]Resultln[BLOCK_SIZE*ARRAY_SIZE-1:0],
	input [3:0]mask[ARRAY_SIZE*ARRAY_SIZE-1:0],
	input Block_control,
	input Direction,
	input Control,
	input ResultCapture,
	input Clk,
	input rst,
	output [4*DATA_WIDTH-1:0]Array_Output[BLOCK_SIZE*ARRAY_SIZE-1:0]
	);
	
	wire [4*DATA_WIDTH-1:0]Array_process[4*(BLOCK_SIZE-1)*BLOCK_SIZE-1:0];
	
	
	//The first column
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_00
	(
		.Input_act_data(Input_act[0]),
		.Input_weight(Input_weight[0]),
		.mask(mask[0]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Resultln[0]),
		.ResultIn_1(Resultln[1]),
		.ResultIn_2(Resultln[2]),
		.ResultIn_2(Resultln[3]),
		.Cell_Output_data_0(Array_process[0]),
		.Cell_Output_data_1(Array_process[1]),
		.Cell_Output_data_2(Array_process[2]),
		.Cell_Output_data_3(Array_process[3])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_10
	(
		.Input_act_data(Input_act[1]),
		.Input_weight(Input_weight[0]),
		.mask(mask[4]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[0]),
		.ResultIn_1(Array_process[1]),
		.ResultIn_2(Array_process[2]),
		.ResultIn_2(Array_process[3]),
		.Cell_Output_data_0(Array_process[16]),
		.Cell_Output_data_1(Array_process[17]),
		.Cell_Output_data_2(Array_process[18]),
		.Cell_Output_data_3(Array_process[19])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_20
	(
		.Input_act_data(Input_act[2]),
		.Input_weight(Input_weight[0]),
		.mask(mask[8]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[16]),
		.ResultIn_1(Array_process[17]),
		.ResultIn_2(Array_process[18]),
		.ResultIn_2(Array_process[19]),
		.Cell_Output_data_0(Array_process[32]),
		.Cell_Output_data_1(Array_process[33]),
		.Cell_Output_data_2(Array_process[34]),
		.Cell_Output_data_3(Array_process[35])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_30
	(
		.Input_act_data(Input_act[3]),
		.Input_weight(Input_weight[0]),
		.mask(mask[12]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[32]),
		.ResultIn_1(Array_process[33]),
		.ResultIn_2(Array_process[34]),
		.ResultIn_2(Array_process[35]),
		.Cell_Output_data_0(Array_Output[0]),
		.Cell_Output_data_1(Array_Output[1]),
		.Cell_Output_data_2(Array_Output[2]),
		.Cell_Output_data_3(Array_Output[3])
	);
  
	//the second column
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_01
	(
		.Input_act_data(Input_act[0]),
		.Input_weight(Input_weight[1]),
		.mask(mask[1]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Resultln[4]),
		.ResultIn_1(Resultln[5]),
		.ResultIn_2(Resultln[6]),
		.ResultIn_2(Resultln[7]),
		.Cell_Output_data_0(Array_process[4]),
		.Cell_Output_data_1(Array_process[5]),
		.Cell_Output_data_2(Array_process[6]),
		.Cell_Output_data_3(Array_process[7])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_11
	(
		.Input_act_data(Input_act[1]),
		.Input_weight(Input_weight[1]),
		.mask(mask[5]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[4]),
		.ResultIn_1(Array_process[5]),
		.ResultIn_2(Array_process[6]),
		.ResultIn_2(Array_process[7]),
		.Cell_Output_data_0(Array_process[20]),
		.Cell_Output_data_1(Array_process[21]),
		.Cell_Output_data_2(Array_process[22]),
		.Cell_Output_data_3(Array_process[23])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_21
	(
		.Input_act_data(Input_act[2]),
		.Input_weight(Input_weight[1]),
		.mask(mask[9]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[20]),
		.ResultIn_1(Array_process[21]),
		.ResultIn_2(Array_process[22]),
		.ResultIn_2(Array_process[23]),
		.Cell_Output_data_0(Array_process[36]),
		.Cell_Output_data_1(Array_process[37]),
		.Cell_Output_data_2(Array_process[38]),
		.Cell_Output_data_3(Array_process[39])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_31
	(
		.Input_act_data(Input_act[3]),
		.Input_weight(Input_weight[1]),
		.mask(mask[13]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[36]),
		.ResultIn_1(Array_process[37]),
		.ResultIn_2(Array_process[38]),
		.ResultIn_2(Array_process[39]),
		.Cell_Output_data_0(Array_Output[4]),
		.Cell_Output_data_1(Array_Output[5]),
		.Cell_Output_data_2(Array_Output[6]),
		.Cell_Output_data_3(Array_Output[7])
	);
  	
	//the third column
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_02
	(
		.Input_act_data(Input_act[0]),
		.Input_weight(Input_weight[2]),
		.mask(mask[2]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Resultln[8]),
		.ResultIn_1(Resultln[9]),
		.ResultIn_2(Resultln[10]),
		.ResultIn_2(Resultln[11]),
		.Cell_Output_data_0(Array_process[8]),
		.Cell_Output_data_1(Array_process[9]),
		.Cell_Output_data_2(Array_process[10]),
		.Cell_Output_data_3(Array_process[11])
	);

	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_12
	(
		.Input_act_data(Input_act[1]),
		.Input_weight(Input_weight[2]),
		.mask(mask[6]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[8]),
		.ResultIn_1(Array_process[9]),
		.ResultIn_2(Array_process[10]),
		.ResultIn_2(Array_process[11]),
		.Cell_Output_data_0(Array_process[24]),
		.Cell_Output_data_1(Array_process[25]),
		.Cell_Output_data_2(Array_process[26]),
		.Cell_Output_data_3(Array_process[27])
	);
  	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_22
	(
		.Input_act_data(Input_act[2]),
		.Input_weight(Input_weight[2]),
		.mask(mask[10]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[24]),
		.ResultIn_1(Array_process[25]),
		.ResultIn_2(Array_process[26]),
		.ResultIn_2(Array_process[27]),
		.Cell_Output_data_0(Array_process[40]),
		.Cell_Output_data_1(Array_process[41]),
		.Cell_Output_data_2(Array_process[42]),
		.Cell_Output_data_3(Array_process[43])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_32
	(
		.Input_act_data(Input_act[3]),
		.Input_weight(Input_weight[2]),
		.mask(mask[14]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[40]),
		.ResultIn_1(Array_process[41]),
		.ResultIn_2(Array_process[42]),
		.ResultIn_2(Array_process[43]),
		.Cell_Output_data_0(Array_Output[8]),
		.Cell_Output_data_1(Array_Output[9]),
		.Cell_Output_data_2(Array_Output[10]),
		.Cell_Output_data_3(Array_Output[11])
	);
  	
	//the fouth column
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_03
	(
		.Input_act_data(Input_act[0]),
		.Input_weight(Input_weight[3]),
		.mask(mask[3]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Resultln[12]),
		.ResultIn_1(Resultln[13]),
		.ResultIn_2(Resultln[14]),
		.ResultIn_2(Resultln[15]),
		.Cell_Output_data_0(Array_process[12]),
		.Cell_Output_data_1(Array_process[13]),
		.Cell_Output_data_2(Array_process[14]),
		.Cell_Output_data_3(Array_process[15])
	);

	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_13
	(
		.Input_act_data(Input_act[1]),
		.Input_weight(Input_weight[3]),
		.mask(mask[7]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[12]),
		.ResultIn_1(Array_process[13]),
		.ResultIn_2(Array_process[14]),
		.ResultIn_2(Array_process[15]),
		.Cell_Output_data_0(Array_process[28]),
		.Cell_Output_data_1(Array_process[29]),
		.Cell_Output_data_2(Array_process[30]),
		.Cell_Output_data_3(Array_process[31])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_23
	(
		.Input_act_data(Input_act[2]),
		.Input_weight(Input_weight[3]),
		.mask(mask[11]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[18]),
		.ResultIn_1(Array_process[29]),
		.ResultIn_2(Array_process[30]),
		.ResultIn_2(Array_process[31]),
		.Cell_Output_data_0(Array_process[44]),
		.Cell_Output_data_1(Array_process[45]),
		.Cell_Output_data_2(Array_process[46]),
		.Cell_Output_data_3(Array_process[47])
	);
	
	CELL_UNIT
	#(
		.DATA_WIDTH(DATA_WIDTH),
		.BLOCK_SIZE(BLOCK_SIZE),
		.SELECT_WIDTH(SELECT_WIDTH)
	)
	Cell_unit_33
	(
		.Input_act_data(Input_act[3]),
		.Input_weight(Input_weight[3]),
		.mask(mask[15]),
		.Block_control(Block_control),
		.Direction(Direction),
		.Control(Control),
		.ResultCapture(ResultCapture),
		.Clk(Clk),
		.rst(rst),
		.ResultIn_0(Array_process[44]),
		.ResultIn_1(Array_process[45]),
		.ResultIn_2(Array_process[46]),
		.ResultIn_2(Array_process[47]),
		.Cell_Output_data_0(Array_Output[12]),
		.Cell_Output_data_1(Array_Output[13]),
		.Cell_Output_data_2(Array_Output[14]),
		.Cell_Output_data_3(Array_Output[15])
	);
endmodule 
  	
	
